grammar edu:umn:cs:melt:exts:ableC:goConcurrency:src:concretesyntax:arrow;

imports edu:umn:cs:melt:ableC:concretesyntax only Ckeyword;

marking terminal Arrow_t '<-' lexer classes{Ckeyword};