grammar edu:umn:cs:melt:exts:ableC:goConcurrency:concretesyntax;

exports edu:umn:cs:melt:exts:ableC:goConcurrency:concretesyntax:close;
exports edu:umn:cs:melt:exts:ableC:goConcurrency:concretesyntax:send;
exports edu:umn:cs:melt:exts:ableC:goConcurrency:concretesyntax:recieve;
exports edu:umn:cs:melt:exts:ableC:goConcurrency:concretesyntax:spawn;
exports edu:umn:cs:melt:exts:ableC:goConcurrency:concretesyntax:select;