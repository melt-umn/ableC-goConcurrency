grammar edu:umn:cs:melt:exts:ableC:goConcurrency:concretesyntax:selectAssignTerm;

imports edu:umn:cs:melt:ableC:concretesyntax only Ckeyword;

terminal Test_t '<==' lexer classes{Ckeyword};