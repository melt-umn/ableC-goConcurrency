grammar edu:umn:cs:melt:exts:ableC:goConcurrency:concretesyntax:closeTerm;

imports edu:umn:cs:melt:ableC:concretesyntax only Ckeyword;

marking terminal Close_t 'close' lexer classes {Ckeyword};