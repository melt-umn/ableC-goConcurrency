grammar determinism;

import edu:umn:cs:melt:ableC:host ;

copper_mda testRecieve(ablecParser) {
  edu:umn:cs:melt:exts:ableC:goConcurrency:concretesyntax:channel;
}

copper_mda testSpawn(ablecParser) {
  edu:umn:cs:melt:exts:ableC:goConcurrency:concretesyntax:spawn;
}