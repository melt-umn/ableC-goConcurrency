grammar edu:umn:cs:melt:exts:ableC:goConcurrency;

exports edu:umn:cs:melt:exts:ableC:goConcurrency:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:goConcurrency:concretesyntax;