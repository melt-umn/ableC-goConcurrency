grammar edu:umn:cs:melt:exts:ableC:goConcurrency:src;

exports edu:umn:cs:melt:exts:ableC:goConcurrency:src:abstractsyntax;

exports edu:umn:cs:melt:exts:ableC:goConcurrency:src:concretesyntax:arrow;
exports edu:umn:cs:melt:exts:ableC:goConcurrency:src:concretesyntax:arrowInfix;
exports edu:umn:cs:melt:exts:ableC:goConcurrency:src:concretesyntax:closeTerm;
exports edu:umn:cs:melt:exts:ableC:goConcurrency:src:concretesyntax:close;
exports edu:umn:cs:melt:exts:ableC:goConcurrency:src:concretesyntax:send;
exports edu:umn:cs:melt:exts:ableC:goConcurrency:src:concretesyntax:recieve;
exports edu:umn:cs:melt:exts:ableC:goConcurrency:src:concretesyntax:spawnTerm;
exports edu:umn:cs:melt:exts:ableC:goConcurrency:src:concretesyntax:spawn;
exports edu:umn:cs:melt:exts:ableC:goConcurrency:src:concretesyntax:selectCases;
exports edu:umn:cs:melt:exts:ableC:goConcurrency:src:concretesyntax:selectExpr;
exports edu:umn:cs:melt:exts:ableC:goConcurrency:src:concretesyntax:selectAssignTerm;
exports edu:umn:cs:melt:exts:ableC:goConcurrency:src:concretesyntax:selectTerm;
exports edu:umn:cs:melt:exts:ableC:goConcurrency:src:concretesyntax:select;
