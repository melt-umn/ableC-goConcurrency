grammar edu:umn:cs:melt:exts:ableC:goConcurrency:src:abstractsyntax;

imports silver:langutil:pp;

nonterminal SelectExpr with location, pp, value, chanType, chan;
nonterminal SelectCases with location, pp, errors, body, lifted<SelectCases>, globalDecls, env, def;

synthesized attribute value::Expr;
synthesized attribute chan::Expr;
synthesized attribute chanType::String;
synthesized attribute body::Stmt;
synthesized attribute def::Maybe<Stmt>;

abstract production chanCond 
top::Expr ::= chExpr::SelectExpr 
{
  forwards to if chExpr.chanType == "receive" then tryReceive(chExpr.chan, location=top.location)
    else if chExpr.chanType == "send" then trySend(chExpr.chan, chExpr.value, location=top.location)
     else tryAssign(chExpr.chan, chExpr.value, location=top.location);
}

abstract production makeReceive
top::SelectExpr ::= ch::Expr
{
  top.chanType = "receive";
  top.chan = ch;
  top.value = ch;
  top.pp = text("receive");
}

abstract production makeSend
top::SelectExpr ::= ch::Expr v::Expr
{
  top.chanType = "send";
  top.chan = ch;
  top.value = v;
  top.pp = text("send");
}

abstract production makeAssign
top::SelectExpr ::= ch::Expr v::Expr
{
  top.chanType = "assign";
  top.chan = ch;
  top.value = v;
  top.pp = text("assign");
}

abstract production trySend
top::Expr ::= ch::Expr v::Expr
{
  forwards to 
      callExpr(
          tmp:templateDeclRefExpr(name("chan_send_select",location=top.location), 
              consTypeName(typeName(directTypeExpr(v.typerep), baseTypeExpr()),
                   nilTypeName()),location=top.location),
          consExpr(ch, consExpr(v, nilExpr())), location=top.location);
}

abstract production tryAssign
top::Expr ::= ch::Expr v::Expr
{
  local channelType::Type = channelSubType(ch.typerep, ch.env);

  forwards to 
      callExpr(
          tmp:templateDeclRefExpr(name("chan_recv_select",location=top.location), 
              consTypeName(typeName(directTypeExpr(channelType), baseTypeExpr()),
                   nilTypeName()),location=top.location),
                                               -- this v needs to be the pointer to v!
          consExpr(ch, consExpr(v, nilExpr())), location=top.location);
}

abstract production tryReceive
top::Expr ::= ch::Expr
{
  local channelType::Type = channelSubType(ch.typerep, ch.env);

  forwards to 
      callExpr(
          tmp:templateDeclRefExpr(name("chan_recv_select_drop",location=top.location), 
              consTypeName(typeName(directTypeExpr(channelType), baseTypeExpr()),
                   nilTypeName()),location=top.location),
          consExpr(ch, nilExpr()), location=top.location);
}

abstract production select
top::Stmt ::= cs::SelectCases {
  
   local body::Stmt = case cs.def of 
                 just(def) -> seqStmt(cs.body, def) 
               | nothing() -> cs.body end;
     
   forwards to whileStmt(
            mkIntConst(1, cs.location),
            body);  
}


abstract production nilCase
top::SelectCases ::= {
   propagate lifted;
   top.pp = text("");
   top.errors := [];
   top.globalDecls := [];
   top.def = nothing();
   top.body = nullStmt();
}

abstract production chanCase 
top::SelectCases ::= chexp::SelectExpr stm::Stmt sc::SelectCases {
   propagate lifted;
   top.globalDecls := sc.globalDecls;
   top.def = sc.def;
   top.pp = ppConcat([chexp.pp, sc.pp]);
   top.errors := sc.errors;

   sc.env = top.env;
   top.body = seqStmt(
                ifStmtNoElse(
                        chanCond(chexp, location=top.location),
                        seqStmt(stm,breakStmt())),
                sc.body);
}

abstract production defaultCase 
top::SelectCases ::= stm::Stmt sc::SelectCases {
   propagate lifted;
   top.body = sc.body;
   top.pp = ppConcat([text("default,"), sc.pp]);

   top.def = case sc.def of 
       just(def) -> nothing()
     | nothing() -> just(seqStmt(stm, breakStmt())) end;
   
   top.errors := sc.errors;
   --top.errors <- case top.def of
   --  nothing() then "Multiple default statements in select" ++ top.errors
   --             else top.errors;
}