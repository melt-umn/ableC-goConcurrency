grammar edu:umn:cs:melt:exts:ableC:goConcurrency:src:concretesyntax:arrowInfix;

imports edu:umn:cs:melt:exts:ableC:goConcurrency:src:concretesyntax:arrow;

nonterminal ArrowInfix_c;

concrete production arrowInfix
top::ArrowInfix_c ::= '<-' 
{
} 