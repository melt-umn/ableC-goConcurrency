grammar edu:umn:cs:melt:exts:ableC:goConcurrency:concretesyntax;

exports edu:umn:cs:melt:exts:ableC:goConcurrency:concretesyntax:channel;
exports edu:umn:cs:melt:exts:ableC:goConcurrency:concretesyntax:spawn;