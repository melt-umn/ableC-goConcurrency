grammar edu:umn:cs:melt:exts:ableC:goConcurrency:concretesyntax:arrowInfix;

exports edu:umn:cs:melt:exts:ableC:goConcurrency:concretesyntax:arrow;

nonterminal ArrowInfix_c;

concrete production arrowInfix
top::ArrowInfix_c ::= '<-' 
{
} 