grammar edu:umn:cs:melt:exts:ableC:goConcurrency:src ;

exports edu:umn:cs:melt:exts:ableC:goConcurrency:src:abstractsyntax ;
exports edu:umn:cs:melt:exts:ableC:goConcurrency:src:concretesyntax ;

