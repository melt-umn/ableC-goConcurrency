grammar edu:umn:cs:melt:exts:ableC:goConcurrency:concretesyntax:selectTerm;

imports edu:umn:cs:melt:ableC:concretesyntax only Ckeyword;

marking terminal Select_t 'select' lexer classes{Ckeyword};