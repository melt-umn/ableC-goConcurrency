grammar edu:umn:cs:melt:exts:ableC:goConcurrency:src:concretesyntax:spawnTerm;

imports edu:umn:cs:melt:ableC:concretesyntax only Ckeyword;

marking terminal Spawn_t 'spawn' lexer classes {Ckeyword};