grammar edu:umn:cs:melt:exts:ableC:goConcurrency:concretesyntax:arrow;

imports edu:umn:cs:melt:ableC:concretesyntax only Cassignment;

marking terminal Arrow_t '<-' lexer classes{Cassignment }, association = left;