grammar edu:umn:cs:melt:exts:ableC:goConcurrency:src ;

exports edu:umn:cs:melt:exts:ableC:goConcurrency:src:abstractsyntax;

exports edu:umn:cs:melt:exts:ableC:goConcurrency:src:concretesyntax:arrow;
exports edu:umn:cs:melt:exts:ableC:goConcurrency:src:concretesyntax:channel;
exports edu:umn:cs:melt:exts:ableC:goConcurrency:src:concretesyntax:spawn;
exports edu:umn:cs:melt:exts:ableC:goConcurrency:src:concretesyntax:select;